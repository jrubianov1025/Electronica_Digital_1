module TOP_Multiplicador (

    input reset,
    input clk,
    input init,

    input [15:0] Multiplicando,
    input [15:0] Multiplicador,
    
    output [31:0] Resultado,
    output DONE

);

wire W_LD;
wire W_SH;
wire W_ADD;
wire W_DEC;
wire W_Z;
wire W_LSB;





endmodule
